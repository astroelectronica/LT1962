.title KiCad schematic
.include "C:/AE/LT1962/_models/C3216X5R2A105K160AA_s.mod"
.include "C:/AE/LT1962/_models/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/LT1962/_models/CGA5L3X5R1H106K160AB_s.mod"
.include "C:/AE/LT1962/_models/LT1962.lib"
R2 /VOUT /ADJ {RADJU}
R3 /ADJ 0 {RADJB}
I1 /VOUT 0 {ILOAD}
XU3 /VOUT 0 CGA5L3X5R1H106K160AB_s
XU4 /BYP /VOUT CEU4J2X7R2A103K125AE_s
V1 /VIN 0 {VSOURCE}
XU1 /VIN 0 C3216X5R2A105K160AA_s
XU2 /VOUT /ADJ /BYP 0 /VIN /VIN LT1962
.end
